// final_project.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module final_project (
		input  wire        accumulate_wire_export,         //         accumulate_wire.export
		input  wire        clk_clk,                        //                     clk.clk
		output wire [15:0] grid_pio0_export,               //               grid_pio0.export
		output wire [15:0] grid_pio1_export,               //               grid_pio1.export
		output wire [15:0] grid_pio10_export,              //              grid_pio10.export
		output wire [15:0] grid_pio11_export,              //              grid_pio11.export
		output wire [15:0] grid_pio12_export,              //              grid_pio12.export
		output wire [15:0] grid_pio13_export,              //              grid_pio13.export
		output wire [15:0] grid_pio14_export,              //              grid_pio14.export
		output wire [15:0] grid_pio15_export,              //              grid_pio15.export
		output wire [15:0] grid_pio2_export,               //               grid_pio2.export
		output wire [15:0] grid_pio3_export,               //               grid_pio3.export
		output wire [15:0] grid_pio4_export,               //               grid_pio4.export
		output wire [15:0] grid_pio5_export,               //               grid_pio5.export
		output wire [15:0] grid_pio6_export,               //               grid_pio6.export
		output wire [15:0] grid_pio7_export,               //               grid_pio7.export
		output wire [15:0] grid_pio8_export,               //               grid_pio8.export
		output wire [15:0] grid_pio9_export,               //               grid_pio9.export
		output wire [15:0] hex_digits_export,              //              hex_digits.export
		input  wire [1:0]  key_external_connection_export, // key_external_connection.export
		output wire [7:0]  keycode_export,                 //                 keycode.export
		output wire [13:0] leds_export,                    //                    leds.export
		input  wire        reset_reset_n,                  //                   reset.reset_n
		output wire        sdram_clk_clk,                  //               sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                //              sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                  //                        .ba
		output wire        sdram_wire_cas_n,               //                        .cas_n
		output wire        sdram_wire_cke,                 //                        .cke
		output wire        sdram_wire_cs_n,                //                        .cs_n
		inout  wire [15:0] sdram_wire_dq,                  //                        .dq
		output wire [1:0]  sdram_wire_dqm,                 //                        .dqm
		output wire        sdram_wire_ras_n,               //                        .ras_n
		output wire        sdram_wire_we_n,                //                        .we_n
		input  wire        spi0_MISO,                      //                    spi0.MISO
		output wire        spi0_MOSI,                      //                        .MOSI
		output wire        spi0_SCLK,                      //                        .SCLK
		output wire        spi0_SS_n,                      //                        .SS_n
		input  wire        usb_gpx_export,                 //                 usb_gpx.export
		input  wire        usb_irq_export,                 //                 usb_irq.export
		output wire        usb_rst_export,                 //                 usb_rst.export
		output wire [1:0]  win_pio_export                  //                 win_pio.export
	);

	wire         sdram_pll_c0_clk;                                           // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;      // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;       // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;             // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;              // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                 // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;            // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;           // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;              // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;           // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;            // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_accumulate_s1_readdata;                   // accumulate:readdata -> mm_interconnect_0:accumulate_s1_readdata
	wire   [1:0] mm_interconnect_0_accumulate_s1_address;                    // mm_interconnect_0:accumulate_s1_address -> accumulate:address
	wire         mm_interconnect_0_keycode_s1_chipselect;                    // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                      // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                       // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                         // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                     // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire  [31:0] mm_interconnect_0_usb_irq_s1_readdata;                      // usb_irq:readdata -> mm_interconnect_0:usb_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_irq_s1_address;                       // mm_interconnect_0:usb_irq_s1_address -> usb_irq:address
	wire  [31:0] mm_interconnect_0_usb_gpx_s1_readdata;                      // usb_gpx:readdata -> mm_interconnect_0:usb_gpx_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_gpx_s1_address;                       // mm_interconnect_0:usb_gpx_s1_address -> usb_gpx:address
	wire         mm_interconnect_0_usb_rst_s1_chipselect;                    // mm_interconnect_0:usb_rst_s1_chipselect -> usb_rst:chipselect
	wire  [31:0] mm_interconnect_0_usb_rst_s1_readdata;                      // usb_rst:readdata -> mm_interconnect_0:usb_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_rst_s1_address;                       // mm_interconnect_0:usb_rst_s1_address -> usb_rst:address
	wire         mm_interconnect_0_usb_rst_s1_write;                         // mm_interconnect_0:usb_rst_s1_write -> usb_rst:write_n
	wire  [31:0] mm_interconnect_0_usb_rst_s1_writedata;                     // mm_interconnect_0:usb_rst_s1_writedata -> usb_rst:writedata
	wire         mm_interconnect_0_hex_digits_pio_s1_chipselect;             // mm_interconnect_0:hex_digits_pio_s1_chipselect -> hex_digits_pio:chipselect
	wire  [31:0] mm_interconnect_0_hex_digits_pio_s1_readdata;               // hex_digits_pio:readdata -> mm_interconnect_0:hex_digits_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_digits_pio_s1_address;                // mm_interconnect_0:hex_digits_pio_s1_address -> hex_digits_pio:address
	wire         mm_interconnect_0_hex_digits_pio_s1_write;                  // mm_interconnect_0:hex_digits_pio_s1_write -> hex_digits_pio:write_n
	wire  [31:0] mm_interconnect_0_hex_digits_pio_s1_writedata;              // mm_interconnect_0:hex_digits_pio_s1_writedata -> hex_digits_pio:writedata
	wire         mm_interconnect_0_leds_pio_s1_chipselect;                   // mm_interconnect_0:leds_pio_s1_chipselect -> leds_pio:chipselect
	wire  [31:0] mm_interconnect_0_leds_pio_s1_readdata;                     // leds_pio:readdata -> mm_interconnect_0:leds_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_pio_s1_address;                      // mm_interconnect_0:leds_pio_s1_address -> leds_pio:address
	wire         mm_interconnect_0_leds_pio_s1_write;                        // mm_interconnect_0:leds_pio_s1_write -> leds_pio:write_n
	wire  [31:0] mm_interconnect_0_leds_pio_s1_writedata;                    // mm_interconnect_0:leds_pio_s1_writedata -> leds_pio:writedata
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                          // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                           // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_timer_s1_chipselect;                      // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                        // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_s1_address;                         // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                           // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                       // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_grid_pio0_s1_chipselect;                  // mm_interconnect_0:grid_pio0_s1_chipselect -> grid_pio0:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio0_s1_readdata;                    // grid_pio0:readdata -> mm_interconnect_0:grid_pio0_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio0_s1_address;                     // mm_interconnect_0:grid_pio0_s1_address -> grid_pio0:address
	wire         mm_interconnect_0_grid_pio0_s1_write;                       // mm_interconnect_0:grid_pio0_s1_write -> grid_pio0:write_n
	wire  [31:0] mm_interconnect_0_grid_pio0_s1_writedata;                   // mm_interconnect_0:grid_pio0_s1_writedata -> grid_pio0:writedata
	wire         mm_interconnect_0_grid_pio1_s1_chipselect;                  // mm_interconnect_0:grid_pio1_s1_chipselect -> grid_pio1:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio1_s1_readdata;                    // grid_pio1:readdata -> mm_interconnect_0:grid_pio1_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio1_s1_address;                     // mm_interconnect_0:grid_pio1_s1_address -> grid_pio1:address
	wire         mm_interconnect_0_grid_pio1_s1_write;                       // mm_interconnect_0:grid_pio1_s1_write -> grid_pio1:write_n
	wire  [31:0] mm_interconnect_0_grid_pio1_s1_writedata;                   // mm_interconnect_0:grid_pio1_s1_writedata -> grid_pio1:writedata
	wire         mm_interconnect_0_grid_pio2_s1_chipselect;                  // mm_interconnect_0:grid_pio2_s1_chipselect -> grid_pio2:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio2_s1_readdata;                    // grid_pio2:readdata -> mm_interconnect_0:grid_pio2_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio2_s1_address;                     // mm_interconnect_0:grid_pio2_s1_address -> grid_pio2:address
	wire         mm_interconnect_0_grid_pio2_s1_write;                       // mm_interconnect_0:grid_pio2_s1_write -> grid_pio2:write_n
	wire  [31:0] mm_interconnect_0_grid_pio2_s1_writedata;                   // mm_interconnect_0:grid_pio2_s1_writedata -> grid_pio2:writedata
	wire         mm_interconnect_0_grid_pio3_s1_chipselect;                  // mm_interconnect_0:grid_pio3_s1_chipselect -> grid_pio3:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio3_s1_readdata;                    // grid_pio3:readdata -> mm_interconnect_0:grid_pio3_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio3_s1_address;                     // mm_interconnect_0:grid_pio3_s1_address -> grid_pio3:address
	wire         mm_interconnect_0_grid_pio3_s1_write;                       // mm_interconnect_0:grid_pio3_s1_write -> grid_pio3:write_n
	wire  [31:0] mm_interconnect_0_grid_pio3_s1_writedata;                   // mm_interconnect_0:grid_pio3_s1_writedata -> grid_pio3:writedata
	wire         mm_interconnect_0_grid_pio4_s1_chipselect;                  // mm_interconnect_0:grid_pio4_s1_chipselect -> grid_pio4:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio4_s1_readdata;                    // grid_pio4:readdata -> mm_interconnect_0:grid_pio4_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio4_s1_address;                     // mm_interconnect_0:grid_pio4_s1_address -> grid_pio4:address
	wire         mm_interconnect_0_grid_pio4_s1_write;                       // mm_interconnect_0:grid_pio4_s1_write -> grid_pio4:write_n
	wire  [31:0] mm_interconnect_0_grid_pio4_s1_writedata;                   // mm_interconnect_0:grid_pio4_s1_writedata -> grid_pio4:writedata
	wire         mm_interconnect_0_grid_pio5_s1_chipselect;                  // mm_interconnect_0:grid_pio5_s1_chipselect -> grid_pio5:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio5_s1_readdata;                    // grid_pio5:readdata -> mm_interconnect_0:grid_pio5_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio5_s1_address;                     // mm_interconnect_0:grid_pio5_s1_address -> grid_pio5:address
	wire         mm_interconnect_0_grid_pio5_s1_write;                       // mm_interconnect_0:grid_pio5_s1_write -> grid_pio5:write_n
	wire  [31:0] mm_interconnect_0_grid_pio5_s1_writedata;                   // mm_interconnect_0:grid_pio5_s1_writedata -> grid_pio5:writedata
	wire         mm_interconnect_0_grid_pio6_s1_chipselect;                  // mm_interconnect_0:grid_pio6_s1_chipselect -> grid_pio6:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio6_s1_readdata;                    // grid_pio6:readdata -> mm_interconnect_0:grid_pio6_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio6_s1_address;                     // mm_interconnect_0:grid_pio6_s1_address -> grid_pio6:address
	wire         mm_interconnect_0_grid_pio6_s1_write;                       // mm_interconnect_0:grid_pio6_s1_write -> grid_pio6:write_n
	wire  [31:0] mm_interconnect_0_grid_pio6_s1_writedata;                   // mm_interconnect_0:grid_pio6_s1_writedata -> grid_pio6:writedata
	wire         mm_interconnect_0_grid_pio7_s1_chipselect;                  // mm_interconnect_0:grid_pio7_s1_chipselect -> grid_pio7:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio7_s1_readdata;                    // grid_pio7:readdata -> mm_interconnect_0:grid_pio7_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio7_s1_address;                     // mm_interconnect_0:grid_pio7_s1_address -> grid_pio7:address
	wire         mm_interconnect_0_grid_pio7_s1_write;                       // mm_interconnect_0:grid_pio7_s1_write -> grid_pio7:write_n
	wire  [31:0] mm_interconnect_0_grid_pio7_s1_writedata;                   // mm_interconnect_0:grid_pio7_s1_writedata -> grid_pio7:writedata
	wire         mm_interconnect_0_grid_pio8_s1_chipselect;                  // mm_interconnect_0:grid_pio8_s1_chipselect -> grid_pio8:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio8_s1_readdata;                    // grid_pio8:readdata -> mm_interconnect_0:grid_pio8_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio8_s1_address;                     // mm_interconnect_0:grid_pio8_s1_address -> grid_pio8:address
	wire         mm_interconnect_0_grid_pio8_s1_write;                       // mm_interconnect_0:grid_pio8_s1_write -> grid_pio8:write_n
	wire  [31:0] mm_interconnect_0_grid_pio8_s1_writedata;                   // mm_interconnect_0:grid_pio8_s1_writedata -> grid_pio8:writedata
	wire         mm_interconnect_0_grid_pio9_s1_chipselect;                  // mm_interconnect_0:grid_pio9_s1_chipselect -> grid_pio9:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio9_s1_readdata;                    // grid_pio9:readdata -> mm_interconnect_0:grid_pio9_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio9_s1_address;                     // mm_interconnect_0:grid_pio9_s1_address -> grid_pio9:address
	wire         mm_interconnect_0_grid_pio9_s1_write;                       // mm_interconnect_0:grid_pio9_s1_write -> grid_pio9:write_n
	wire  [31:0] mm_interconnect_0_grid_pio9_s1_writedata;                   // mm_interconnect_0:grid_pio9_s1_writedata -> grid_pio9:writedata
	wire         mm_interconnect_0_grid_pio10_s1_chipselect;                 // mm_interconnect_0:grid_pio10_s1_chipselect -> grid_pio10:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio10_s1_readdata;                   // grid_pio10:readdata -> mm_interconnect_0:grid_pio10_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio10_s1_address;                    // mm_interconnect_0:grid_pio10_s1_address -> grid_pio10:address
	wire         mm_interconnect_0_grid_pio10_s1_write;                      // mm_interconnect_0:grid_pio10_s1_write -> grid_pio10:write_n
	wire  [31:0] mm_interconnect_0_grid_pio10_s1_writedata;                  // mm_interconnect_0:grid_pio10_s1_writedata -> grid_pio10:writedata
	wire         mm_interconnect_0_grid_pio11_s1_chipselect;                 // mm_interconnect_0:grid_pio11_s1_chipselect -> grid_pio11:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio11_s1_readdata;                   // grid_pio11:readdata -> mm_interconnect_0:grid_pio11_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio11_s1_address;                    // mm_interconnect_0:grid_pio11_s1_address -> grid_pio11:address
	wire         mm_interconnect_0_grid_pio11_s1_write;                      // mm_interconnect_0:grid_pio11_s1_write -> grid_pio11:write_n
	wire  [31:0] mm_interconnect_0_grid_pio11_s1_writedata;                  // mm_interconnect_0:grid_pio11_s1_writedata -> grid_pio11:writedata
	wire         mm_interconnect_0_grid_pio12_s1_chipselect;                 // mm_interconnect_0:grid_pio12_s1_chipselect -> grid_pio12:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio12_s1_readdata;                   // grid_pio12:readdata -> mm_interconnect_0:grid_pio12_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio12_s1_address;                    // mm_interconnect_0:grid_pio12_s1_address -> grid_pio12:address
	wire         mm_interconnect_0_grid_pio12_s1_write;                      // mm_interconnect_0:grid_pio12_s1_write -> grid_pio12:write_n
	wire  [31:0] mm_interconnect_0_grid_pio12_s1_writedata;                  // mm_interconnect_0:grid_pio12_s1_writedata -> grid_pio12:writedata
	wire         mm_interconnect_0_grid_pio13_s1_chipselect;                 // mm_interconnect_0:grid_pio13_s1_chipselect -> grid_pio13:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio13_s1_readdata;                   // grid_pio13:readdata -> mm_interconnect_0:grid_pio13_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio13_s1_address;                    // mm_interconnect_0:grid_pio13_s1_address -> grid_pio13:address
	wire         mm_interconnect_0_grid_pio13_s1_write;                      // mm_interconnect_0:grid_pio13_s1_write -> grid_pio13:write_n
	wire  [31:0] mm_interconnect_0_grid_pio13_s1_writedata;                  // mm_interconnect_0:grid_pio13_s1_writedata -> grid_pio13:writedata
	wire         mm_interconnect_0_grid_pio14_s1_chipselect;                 // mm_interconnect_0:grid_pio14_s1_chipselect -> grid_pio14:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio14_s1_readdata;                   // grid_pio14:readdata -> mm_interconnect_0:grid_pio14_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio14_s1_address;                    // mm_interconnect_0:grid_pio14_s1_address -> grid_pio14:address
	wire         mm_interconnect_0_grid_pio14_s1_write;                      // mm_interconnect_0:grid_pio14_s1_write -> grid_pio14:write_n
	wire  [31:0] mm_interconnect_0_grid_pio14_s1_writedata;                  // mm_interconnect_0:grid_pio14_s1_writedata -> grid_pio14:writedata
	wire         mm_interconnect_0_grid_pio15_s1_chipselect;                 // mm_interconnect_0:grid_pio15_s1_chipselect -> grid_pio15:chipselect
	wire  [31:0] mm_interconnect_0_grid_pio15_s1_readdata;                   // grid_pio15:readdata -> mm_interconnect_0:grid_pio15_s1_readdata
	wire   [1:0] mm_interconnect_0_grid_pio15_s1_address;                    // mm_interconnect_0:grid_pio15_s1_address -> grid_pio15:address
	wire         mm_interconnect_0_grid_pio15_s1_write;                      // mm_interconnect_0:grid_pio15_s1_write -> grid_pio15:write_n
	wire  [31:0] mm_interconnect_0_grid_pio15_s1_writedata;                  // mm_interconnect_0:grid_pio15_s1_writedata -> grid_pio15:writedata
	wire         mm_interconnect_0_win_lose_pio_s1_chipselect;               // mm_interconnect_0:win_lose_pio_s1_chipselect -> win_lose_pio:chipselect
	wire  [31:0] mm_interconnect_0_win_lose_pio_s1_readdata;                 // win_lose_pio:readdata -> mm_interconnect_0:win_lose_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_win_lose_pio_s1_address;                  // mm_interconnect_0:win_lose_pio_s1_address -> win_lose_pio:address
	wire         mm_interconnect_0_win_lose_pio_s1_write;                    // mm_interconnect_0:win_lose_pio_s1_write -> win_lose_pio:write_n
	wire  [31:0] mm_interconnect_0_win_lose_pio_s1_writedata;                // mm_interconnect_0:win_lose_pio_s1_writedata -> win_lose_pio:writedata
	wire         mm_interconnect_0_spi0_spi_control_port_chipselect;         // mm_interconnect_0:spi0_spi_control_port_chipselect -> spi0:spi_select
	wire  [15:0] mm_interconnect_0_spi0_spi_control_port_readdata;           // spi0:data_to_cpu -> mm_interconnect_0:spi0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi0_spi_control_port_address;            // mm_interconnect_0:spi0_spi_control_port_address -> spi0:mem_addr
	wire         mm_interconnect_0_spi0_spi_control_port_read;               // mm_interconnect_0:spi0_spi_control_port_read -> spi0:read_n
	wire         mm_interconnect_0_spi0_spi_control_port_write;              // mm_interconnect_0:spi0_spi_control_port_write -> spi0:write_n
	wire  [15:0] mm_interconnect_0_spi0_spi_control_port_writedata;          // mm_interconnect_0:spi0_spi_control_port_writedata -> spi0:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // spi0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [accumulate:reset_n, grid_pio0:reset_n, grid_pio10:reset_n, grid_pio11:reset_n, grid_pio12:reset_n, grid_pio13:reset_n, grid_pio14:reset_n, grid_pio15:reset_n, grid_pio1:reset_n, grid_pio2:reset_n, grid_pio3:reset_n, grid_pio4:reset_n, grid_pio5:reset_n, grid_pio6:reset_n, grid_pio7:reset_n, grid_pio8:reset_n, grid_pio9:reset_n, hex_digits_pio:reset_n, irq_mapper:reset, jtag_uart:rst_n, key:reset_n, keycode:reset_n, leds_pio:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram_pll:reset, spi0:reset_n, sysid_qsys_0:reset_n, timer:reset_n, usb_gpx:reset_n, usb_irq:reset_n, usb_rst:reset_n, win_lose_pio:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	final_project_accumulate accumulate (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_accumulate_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_accumulate_s1_readdata), //                    .readdata
		.in_port  (accumulate_wire_export)                    // external_connection.export
	);

	final_project_grid_pio0 grid_pio0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio0_s1_readdata),   //                    .readdata
		.out_port   (grid_pio0_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio1 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio1_s1_readdata),   //                    .readdata
		.out_port   (grid_pio1_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio10 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio10_s1_readdata),   //                    .readdata
		.out_port   (grid_pio10_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio11 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio11_s1_readdata),   //                    .readdata
		.out_port   (grid_pio11_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio12 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio12_s1_readdata),   //                    .readdata
		.out_port   (grid_pio12_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio13 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio13_s1_readdata),   //                    .readdata
		.out_port   (grid_pio13_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio14 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio14_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio14_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio14_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio14_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio14_s1_readdata),   //                    .readdata
		.out_port   (grid_pio14_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio15 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio15_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio15_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio15_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio15_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio15_s1_readdata),   //                    .readdata
		.out_port   (grid_pio15_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio2 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio2_s1_readdata),   //                    .readdata
		.out_port   (grid_pio2_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio3 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio3_s1_readdata),   //                    .readdata
		.out_port   (grid_pio3_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio4 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio4_s1_readdata),   //                    .readdata
		.out_port   (grid_pio4_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio5 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio5_s1_readdata),   //                    .readdata
		.out_port   (grid_pio5_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio6 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio6_s1_readdata),   //                    .readdata
		.out_port   (grid_pio6_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio7 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio7_s1_readdata),   //                    .readdata
		.out_port   (grid_pio7_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio8 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio8_s1_readdata),   //                    .readdata
		.out_port   (grid_pio8_export)                           // external_connection.export
	);

	final_project_grid_pio0 grid_pio9 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_grid_pio9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_grid_pio9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_grid_pio9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_grid_pio9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_grid_pio9_s1_readdata),   //                    .readdata
		.out_port   (grid_pio9_export)                           // external_connection.export
	);

	final_project_grid_pio0 hex_digits_pio (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_hex_digits_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_digits_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_digits_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_digits_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_digits_pio_s1_readdata),   //                    .readdata
		.out_port   (hex_digits_export)                               // external_connection.export
	);

	final_project_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	final_project_key key (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata), //                    .readdata
		.in_port  (key_external_connection_export)     // external_connection.export
	);

	final_project_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	final_project_leds_pio leds_pio (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_leds_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_pio_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                               // external_connection.export
	);

	final_project_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	final_project_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	final_project_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_project_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.c2                 (),                                                //           (terminated)
		.c3                 (),                                                //           (terminated)
		.c4                 (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (3'b000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	final_project_spi0 spi0 (
		.clk           (clk_clk),                                            //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                    //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                           //              irq.irq
		.MISO          (spi0_MISO),                                          //         external.export
		.MOSI          (spi0_MOSI),                                          //                 .export
		.SCLK          (spi0_SCLK),                                          //                 .export
		.SS_n          (spi0_SS_n)                                           //                 .export
	);

	final_project_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	final_project_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	final_project_accumulate usb_gpx (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_usb_gpx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_gpx_s1_readdata), //                    .readdata
		.in_port  (usb_gpx_export)                         // external_connection.export
	);

	final_project_accumulate usb_irq (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_usb_irq_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_irq_s1_readdata), //                    .readdata
		.in_port  (usb_irq_export)                         // external_connection.export
	);

	final_project_usb_rst usb_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_usb_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_usb_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_usb_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_usb_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_usb_rst_s1_readdata),   //                    .readdata
		.out_port   (usb_rst_export)                           // external_connection.export
	);

	final_project_win_lose_pio win_lose_pio (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_win_lose_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_win_lose_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_win_lose_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_win_lose_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_win_lose_pio_s1_readdata),   //                    .readdata
		.out_port   (win_pio_export)                                // external_connection.export
	);

	final_project_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                           //                             sdram_pll_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                         //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.accumulate_s1_address                          (mm_interconnect_0_accumulate_s1_address),                    //                            accumulate_s1.address
		.accumulate_s1_readdata                         (mm_interconnect_0_accumulate_s1_readdata),                   //                                         .readdata
		.grid_pio0_s1_address                           (mm_interconnect_0_grid_pio0_s1_address),                     //                             grid_pio0_s1.address
		.grid_pio0_s1_write                             (mm_interconnect_0_grid_pio0_s1_write),                       //                                         .write
		.grid_pio0_s1_readdata                          (mm_interconnect_0_grid_pio0_s1_readdata),                    //                                         .readdata
		.grid_pio0_s1_writedata                         (mm_interconnect_0_grid_pio0_s1_writedata),                   //                                         .writedata
		.grid_pio0_s1_chipselect                        (mm_interconnect_0_grid_pio0_s1_chipselect),                  //                                         .chipselect
		.grid_pio1_s1_address                           (mm_interconnect_0_grid_pio1_s1_address),                     //                             grid_pio1_s1.address
		.grid_pio1_s1_write                             (mm_interconnect_0_grid_pio1_s1_write),                       //                                         .write
		.grid_pio1_s1_readdata                          (mm_interconnect_0_grid_pio1_s1_readdata),                    //                                         .readdata
		.grid_pio1_s1_writedata                         (mm_interconnect_0_grid_pio1_s1_writedata),                   //                                         .writedata
		.grid_pio1_s1_chipselect                        (mm_interconnect_0_grid_pio1_s1_chipselect),                  //                                         .chipselect
		.grid_pio10_s1_address                          (mm_interconnect_0_grid_pio10_s1_address),                    //                            grid_pio10_s1.address
		.grid_pio10_s1_write                            (mm_interconnect_0_grid_pio10_s1_write),                      //                                         .write
		.grid_pio10_s1_readdata                         (mm_interconnect_0_grid_pio10_s1_readdata),                   //                                         .readdata
		.grid_pio10_s1_writedata                        (mm_interconnect_0_grid_pio10_s1_writedata),                  //                                         .writedata
		.grid_pio10_s1_chipselect                       (mm_interconnect_0_grid_pio10_s1_chipselect),                 //                                         .chipselect
		.grid_pio11_s1_address                          (mm_interconnect_0_grid_pio11_s1_address),                    //                            grid_pio11_s1.address
		.grid_pio11_s1_write                            (mm_interconnect_0_grid_pio11_s1_write),                      //                                         .write
		.grid_pio11_s1_readdata                         (mm_interconnect_0_grid_pio11_s1_readdata),                   //                                         .readdata
		.grid_pio11_s1_writedata                        (mm_interconnect_0_grid_pio11_s1_writedata),                  //                                         .writedata
		.grid_pio11_s1_chipselect                       (mm_interconnect_0_grid_pio11_s1_chipselect),                 //                                         .chipselect
		.grid_pio12_s1_address                          (mm_interconnect_0_grid_pio12_s1_address),                    //                            grid_pio12_s1.address
		.grid_pio12_s1_write                            (mm_interconnect_0_grid_pio12_s1_write),                      //                                         .write
		.grid_pio12_s1_readdata                         (mm_interconnect_0_grid_pio12_s1_readdata),                   //                                         .readdata
		.grid_pio12_s1_writedata                        (mm_interconnect_0_grid_pio12_s1_writedata),                  //                                         .writedata
		.grid_pio12_s1_chipselect                       (mm_interconnect_0_grid_pio12_s1_chipselect),                 //                                         .chipselect
		.grid_pio13_s1_address                          (mm_interconnect_0_grid_pio13_s1_address),                    //                            grid_pio13_s1.address
		.grid_pio13_s1_write                            (mm_interconnect_0_grid_pio13_s1_write),                      //                                         .write
		.grid_pio13_s1_readdata                         (mm_interconnect_0_grid_pio13_s1_readdata),                   //                                         .readdata
		.grid_pio13_s1_writedata                        (mm_interconnect_0_grid_pio13_s1_writedata),                  //                                         .writedata
		.grid_pio13_s1_chipselect                       (mm_interconnect_0_grid_pio13_s1_chipselect),                 //                                         .chipselect
		.grid_pio14_s1_address                          (mm_interconnect_0_grid_pio14_s1_address),                    //                            grid_pio14_s1.address
		.grid_pio14_s1_write                            (mm_interconnect_0_grid_pio14_s1_write),                      //                                         .write
		.grid_pio14_s1_readdata                         (mm_interconnect_0_grid_pio14_s1_readdata),                   //                                         .readdata
		.grid_pio14_s1_writedata                        (mm_interconnect_0_grid_pio14_s1_writedata),                  //                                         .writedata
		.grid_pio14_s1_chipselect                       (mm_interconnect_0_grid_pio14_s1_chipselect),                 //                                         .chipselect
		.grid_pio15_s1_address                          (mm_interconnect_0_grid_pio15_s1_address),                    //                            grid_pio15_s1.address
		.grid_pio15_s1_write                            (mm_interconnect_0_grid_pio15_s1_write),                      //                                         .write
		.grid_pio15_s1_readdata                         (mm_interconnect_0_grid_pio15_s1_readdata),                   //                                         .readdata
		.grid_pio15_s1_writedata                        (mm_interconnect_0_grid_pio15_s1_writedata),                  //                                         .writedata
		.grid_pio15_s1_chipselect                       (mm_interconnect_0_grid_pio15_s1_chipselect),                 //                                         .chipselect
		.grid_pio2_s1_address                           (mm_interconnect_0_grid_pio2_s1_address),                     //                             grid_pio2_s1.address
		.grid_pio2_s1_write                             (mm_interconnect_0_grid_pio2_s1_write),                       //                                         .write
		.grid_pio2_s1_readdata                          (mm_interconnect_0_grid_pio2_s1_readdata),                    //                                         .readdata
		.grid_pio2_s1_writedata                         (mm_interconnect_0_grid_pio2_s1_writedata),                   //                                         .writedata
		.grid_pio2_s1_chipselect                        (mm_interconnect_0_grid_pio2_s1_chipselect),                  //                                         .chipselect
		.grid_pio3_s1_address                           (mm_interconnect_0_grid_pio3_s1_address),                     //                             grid_pio3_s1.address
		.grid_pio3_s1_write                             (mm_interconnect_0_grid_pio3_s1_write),                       //                                         .write
		.grid_pio3_s1_readdata                          (mm_interconnect_0_grid_pio3_s1_readdata),                    //                                         .readdata
		.grid_pio3_s1_writedata                         (mm_interconnect_0_grid_pio3_s1_writedata),                   //                                         .writedata
		.grid_pio3_s1_chipselect                        (mm_interconnect_0_grid_pio3_s1_chipselect),                  //                                         .chipselect
		.grid_pio4_s1_address                           (mm_interconnect_0_grid_pio4_s1_address),                     //                             grid_pio4_s1.address
		.grid_pio4_s1_write                             (mm_interconnect_0_grid_pio4_s1_write),                       //                                         .write
		.grid_pio4_s1_readdata                          (mm_interconnect_0_grid_pio4_s1_readdata),                    //                                         .readdata
		.grid_pio4_s1_writedata                         (mm_interconnect_0_grid_pio4_s1_writedata),                   //                                         .writedata
		.grid_pio4_s1_chipselect                        (mm_interconnect_0_grid_pio4_s1_chipselect),                  //                                         .chipselect
		.grid_pio5_s1_address                           (mm_interconnect_0_grid_pio5_s1_address),                     //                             grid_pio5_s1.address
		.grid_pio5_s1_write                             (mm_interconnect_0_grid_pio5_s1_write),                       //                                         .write
		.grid_pio5_s1_readdata                          (mm_interconnect_0_grid_pio5_s1_readdata),                    //                                         .readdata
		.grid_pio5_s1_writedata                         (mm_interconnect_0_grid_pio5_s1_writedata),                   //                                         .writedata
		.grid_pio5_s1_chipselect                        (mm_interconnect_0_grid_pio5_s1_chipselect),                  //                                         .chipselect
		.grid_pio6_s1_address                           (mm_interconnect_0_grid_pio6_s1_address),                     //                             grid_pio6_s1.address
		.grid_pio6_s1_write                             (mm_interconnect_0_grid_pio6_s1_write),                       //                                         .write
		.grid_pio6_s1_readdata                          (mm_interconnect_0_grid_pio6_s1_readdata),                    //                                         .readdata
		.grid_pio6_s1_writedata                         (mm_interconnect_0_grid_pio6_s1_writedata),                   //                                         .writedata
		.grid_pio6_s1_chipselect                        (mm_interconnect_0_grid_pio6_s1_chipselect),                  //                                         .chipselect
		.grid_pio7_s1_address                           (mm_interconnect_0_grid_pio7_s1_address),                     //                             grid_pio7_s1.address
		.grid_pio7_s1_write                             (mm_interconnect_0_grid_pio7_s1_write),                       //                                         .write
		.grid_pio7_s1_readdata                          (mm_interconnect_0_grid_pio7_s1_readdata),                    //                                         .readdata
		.grid_pio7_s1_writedata                         (mm_interconnect_0_grid_pio7_s1_writedata),                   //                                         .writedata
		.grid_pio7_s1_chipselect                        (mm_interconnect_0_grid_pio7_s1_chipselect),                  //                                         .chipselect
		.grid_pio8_s1_address                           (mm_interconnect_0_grid_pio8_s1_address),                     //                             grid_pio8_s1.address
		.grid_pio8_s1_write                             (mm_interconnect_0_grid_pio8_s1_write),                       //                                         .write
		.grid_pio8_s1_readdata                          (mm_interconnect_0_grid_pio8_s1_readdata),                    //                                         .readdata
		.grid_pio8_s1_writedata                         (mm_interconnect_0_grid_pio8_s1_writedata),                   //                                         .writedata
		.grid_pio8_s1_chipselect                        (mm_interconnect_0_grid_pio8_s1_chipselect),                  //                                         .chipselect
		.grid_pio9_s1_address                           (mm_interconnect_0_grid_pio9_s1_address),                     //                             grid_pio9_s1.address
		.grid_pio9_s1_write                             (mm_interconnect_0_grid_pio9_s1_write),                       //                                         .write
		.grid_pio9_s1_readdata                          (mm_interconnect_0_grid_pio9_s1_readdata),                    //                                         .readdata
		.grid_pio9_s1_writedata                         (mm_interconnect_0_grid_pio9_s1_writedata),                   //                                         .writedata
		.grid_pio9_s1_chipselect                        (mm_interconnect_0_grid_pio9_s1_chipselect),                  //                                         .chipselect
		.hex_digits_pio_s1_address                      (mm_interconnect_0_hex_digits_pio_s1_address),                //                        hex_digits_pio_s1.address
		.hex_digits_pio_s1_write                        (mm_interconnect_0_hex_digits_pio_s1_write),                  //                                         .write
		.hex_digits_pio_s1_readdata                     (mm_interconnect_0_hex_digits_pio_s1_readdata),               //                                         .readdata
		.hex_digits_pio_s1_writedata                    (mm_interconnect_0_hex_digits_pio_s1_writedata),              //                                         .writedata
		.hex_digits_pio_s1_chipselect                   (mm_interconnect_0_hex_digits_pio_s1_chipselect),             //                                         .chipselect
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                         .chipselect
		.key_s1_address                                 (mm_interconnect_0_key_s1_address),                           //                                   key_s1.address
		.key_s1_readdata                                (mm_interconnect_0_key_s1_readdata),                          //                                         .readdata
		.keycode_s1_address                             (mm_interconnect_0_keycode_s1_address),                       //                               keycode_s1.address
		.keycode_s1_write                               (mm_interconnect_0_keycode_s1_write),                         //                                         .write
		.keycode_s1_readdata                            (mm_interconnect_0_keycode_s1_readdata),                      //                                         .readdata
		.keycode_s1_writedata                           (mm_interconnect_0_keycode_s1_writedata),                     //                                         .writedata
		.keycode_s1_chipselect                          (mm_interconnect_0_keycode_s1_chipselect),                    //                                         .chipselect
		.leds_pio_s1_address                            (mm_interconnect_0_leds_pio_s1_address),                      //                              leds_pio_s1.address
		.leds_pio_s1_write                              (mm_interconnect_0_leds_pio_s1_write),                        //                                         .write
		.leds_pio_s1_readdata                           (mm_interconnect_0_leds_pio_s1_readdata),                     //                                         .readdata
		.leds_pio_s1_writedata                          (mm_interconnect_0_leds_pio_s1_writedata),                    //                                         .writedata
		.leds_pio_s1_chipselect                         (mm_interconnect_0_leds_pio_s1_chipselect),                   //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                         .clken
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                         //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                           //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                            //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                        //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                       //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                      //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                     //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                      //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),              //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                 //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),             //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),            //                                         .writedata
		.spi0_spi_control_port_address                  (mm_interconnect_0_spi0_spi_control_port_address),            //                    spi0_spi_control_port.address
		.spi0_spi_control_port_write                    (mm_interconnect_0_spi0_spi_control_port_write),              //                                         .write
		.spi0_spi_control_port_read                     (mm_interconnect_0_spi0_spi_control_port_read),               //                                         .read
		.spi0_spi_control_port_readdata                 (mm_interconnect_0_spi0_spi_control_port_readdata),           //                                         .readdata
		.spi0_spi_control_port_writedata                (mm_interconnect_0_spi0_spi_control_port_writedata),          //                                         .writedata
		.spi0_spi_control_port_chipselect               (mm_interconnect_0_spi0_spi_control_port_chipselect),         //                                         .chipselect
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),       //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),      //                                         .readdata
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                         //                                 timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                           //                                         .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                        //                                         .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                       //                                         .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect),                      //                                         .chipselect
		.usb_gpx_s1_address                             (mm_interconnect_0_usb_gpx_s1_address),                       //                               usb_gpx_s1.address
		.usb_gpx_s1_readdata                            (mm_interconnect_0_usb_gpx_s1_readdata),                      //                                         .readdata
		.usb_irq_s1_address                             (mm_interconnect_0_usb_irq_s1_address),                       //                               usb_irq_s1.address
		.usb_irq_s1_readdata                            (mm_interconnect_0_usb_irq_s1_readdata),                      //                                         .readdata
		.usb_rst_s1_address                             (mm_interconnect_0_usb_rst_s1_address),                       //                               usb_rst_s1.address
		.usb_rst_s1_write                               (mm_interconnect_0_usb_rst_s1_write),                         //                                         .write
		.usb_rst_s1_readdata                            (mm_interconnect_0_usb_rst_s1_readdata),                      //                                         .readdata
		.usb_rst_s1_writedata                           (mm_interconnect_0_usb_rst_s1_writedata),                     //                                         .writedata
		.usb_rst_s1_chipselect                          (mm_interconnect_0_usb_rst_s1_chipselect),                    //                                         .chipselect
		.win_lose_pio_s1_address                        (mm_interconnect_0_win_lose_pio_s1_address),                  //                          win_lose_pio_s1.address
		.win_lose_pio_s1_write                          (mm_interconnect_0_win_lose_pio_s1_write),                    //                                         .write
		.win_lose_pio_s1_readdata                       (mm_interconnect_0_win_lose_pio_s1_readdata),                 //                                         .readdata
		.win_lose_pio_s1_writedata                      (mm_interconnect_0_win_lose_pio_s1_writedata),                //                                         .writedata
		.win_lose_pio_s1_chipselect                     (mm_interconnect_0_win_lose_pio_s1_chipselect)                //                                         .chipselect
	);

	final_project_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
